module mem #(                   // 
    parameter  ADDR_LEN  = 11   // 
) (
    input  clk, rst,
    input  [ADDR_LEN-1:0] addr, // memory address
    output reg [31:0] rd_data,  // data read out
    input  wr_req,
    input  [31:0] wr_data       // data write in
);
localparam MEM_SIZE = 1<<ADDR_LEN;
reg [31:0] ram_cell[768] ;

always @ (posedge clk or posedge rst)
    if(rst)
        rd_data <= 0;
    else
        rd_data <= ram_cell[addr];

always @ (posedge clk)
    if(wr_req) 
        ram_cell[addr] <= wr_data;

initial begin
    // dst matrix C
    ram_cell[       0] = 32'h0;  // 32'h53970897;
    ram_cell[       1] = 32'h0;  // 32'h35c83245;
    ram_cell[       2] = 32'h0;  // 32'h5ba33747;
    ram_cell[       3] = 32'h0;  // 32'h74791417;
    ram_cell[       4] = 32'h0;  // 32'h5b2ff011;
    ram_cell[       5] = 32'h0;  // 32'hfc07ec25;
    ram_cell[       6] = 32'h0;  // 32'hcf2f4474;
    ram_cell[       7] = 32'h0;  // 32'h31428290;
    ram_cell[       8] = 32'h0;  // 32'hc44a889c;
    ram_cell[       9] = 32'h0;  // 32'h0e6b1cbb;
    ram_cell[      10] = 32'h0;  // 32'h00c6258b;
    ram_cell[      11] = 32'h0;  // 32'h027f511c;
    ram_cell[      12] = 32'h0;  // 32'hf4df0ac2;
    ram_cell[      13] = 32'h0;  // 32'h669fc1a5;
    ram_cell[      14] = 32'h0;  // 32'h9a1bb87b;
    ram_cell[      15] = 32'h0;  // 32'h5767f797;
    ram_cell[      16] = 32'h0;  // 32'hcf3dba46;
    ram_cell[      17] = 32'h0;  // 32'h1cea96ec;
    ram_cell[      18] = 32'h0;  // 32'h279d8fcb;
    ram_cell[      19] = 32'h0;  // 32'hcd006d4e;
    ram_cell[      20] = 32'h0;  // 32'h9d20b95f;
    ram_cell[      21] = 32'h0;  // 32'h8896dd2b;
    ram_cell[      22] = 32'h0;  // 32'hfb407f88;
    ram_cell[      23] = 32'h0;  // 32'hf01229f6;
    ram_cell[      24] = 32'h0;  // 32'he4805c50;
    ram_cell[      25] = 32'h0;  // 32'hc2f6136f;
    ram_cell[      26] = 32'h0;  // 32'he288788d;
    ram_cell[      27] = 32'h0;  // 32'h182eec71;
    ram_cell[      28] = 32'h0;  // 32'ha06e6169;
    ram_cell[      29] = 32'h0;  // 32'he6e99066;
    ram_cell[      30] = 32'h0;  // 32'h4fe03753;
    ram_cell[      31] = 32'h0;  // 32'h5bef9bee;
    ram_cell[      32] = 32'h0;  // 32'ha217b92d;
    ram_cell[      33] = 32'h0;  // 32'h02032ba0;
    ram_cell[      34] = 32'h0;  // 32'h3bbab4a0;
    ram_cell[      35] = 32'h0;  // 32'h3a3716fc;
    ram_cell[      36] = 32'h0;  // 32'ha45a23e2;
    ram_cell[      37] = 32'h0;  // 32'hee1f90a6;
    ram_cell[      38] = 32'h0;  // 32'hbb5103a2;
    ram_cell[      39] = 32'h0;  // 32'h29d25394;
    ram_cell[      40] = 32'h0;  // 32'ha997fcce;
    ram_cell[      41] = 32'h0;  // 32'hc0cb7460;
    ram_cell[      42] = 32'h0;  // 32'h5a2c63b5;
    ram_cell[      43] = 32'h0;  // 32'hcf0239d2;
    ram_cell[      44] = 32'h0;  // 32'ha89efb57;
    ram_cell[      45] = 32'h0;  // 32'h004cbeca;
    ram_cell[      46] = 32'h0;  // 32'h223f97b3;
    ram_cell[      47] = 32'h0;  // 32'h767dc3e2;
    ram_cell[      48] = 32'h0;  // 32'hde2af22b;
    ram_cell[      49] = 32'h0;  // 32'h68c8f71d;
    ram_cell[      50] = 32'h0;  // 32'h4d169bb7;
    ram_cell[      51] = 32'h0;  // 32'hf3067ce6;
    ram_cell[      52] = 32'h0;  // 32'hbb76c489;
    ram_cell[      53] = 32'h0;  // 32'hc341197d;
    ram_cell[      54] = 32'h0;  // 32'h9e331197;
    ram_cell[      55] = 32'h0;  // 32'h55b08dfe;
    ram_cell[      56] = 32'h0;  // 32'h60f1868e;
    ram_cell[      57] = 32'h0;  // 32'h3faca500;
    ram_cell[      58] = 32'h0;  // 32'hd227c4e1;
    ram_cell[      59] = 32'h0;  // 32'h31f15c38;
    ram_cell[      60] = 32'h0;  // 32'h8505d25f;
    ram_cell[      61] = 32'h0;  // 32'h5d7af071;
    ram_cell[      62] = 32'h0;  // 32'hf5a79b83;
    ram_cell[      63] = 32'h0;  // 32'hc266547b;
    ram_cell[      64] = 32'h0;  // 32'h41b0c513;
    ram_cell[      65] = 32'h0;  // 32'ha72c2f84;
    ram_cell[      66] = 32'h0;  // 32'h2bdfec89;
    ram_cell[      67] = 32'h0;  // 32'h25ef5a1d;
    ram_cell[      68] = 32'h0;  // 32'h49efae7e;
    ram_cell[      69] = 32'h0;  // 32'ha9c98443;
    ram_cell[      70] = 32'h0;  // 32'h765360fd;
    ram_cell[      71] = 32'h0;  // 32'hd71ae0eb;
    ram_cell[      72] = 32'h0;  // 32'hcdf5c13b;
    ram_cell[      73] = 32'h0;  // 32'h6b08332e;
    ram_cell[      74] = 32'h0;  // 32'h690e9022;
    ram_cell[      75] = 32'h0;  // 32'hfa90a6db;
    ram_cell[      76] = 32'h0;  // 32'hcb4d3945;
    ram_cell[      77] = 32'h0;  // 32'h5f7e69fa;
    ram_cell[      78] = 32'h0;  // 32'hb0133283;
    ram_cell[      79] = 32'h0;  // 32'hed4e4fed;
    ram_cell[      80] = 32'h0;  // 32'h53d5d45b;
    ram_cell[      81] = 32'h0;  // 32'hfcf0842f;
    ram_cell[      82] = 32'h0;  // 32'ha4240ff2;
    ram_cell[      83] = 32'h0;  // 32'h42575b03;
    ram_cell[      84] = 32'h0;  // 32'haa2c5be4;
    ram_cell[      85] = 32'h0;  // 32'h618a22c8;
    ram_cell[      86] = 32'h0;  // 32'h9eb19084;
    ram_cell[      87] = 32'h0;  // 32'h3ff46989;
    ram_cell[      88] = 32'h0;  // 32'h9b666879;
    ram_cell[      89] = 32'h0;  // 32'h17e5cda8;
    ram_cell[      90] = 32'h0;  // 32'h3aad1fe8;
    ram_cell[      91] = 32'h0;  // 32'h523c9a87;
    ram_cell[      92] = 32'h0;  // 32'h3904e5b4;
    ram_cell[      93] = 32'h0;  // 32'hfff2dead;
    ram_cell[      94] = 32'h0;  // 32'h7e691459;
    ram_cell[      95] = 32'h0;  // 32'hd4689dd0;
    ram_cell[      96] = 32'h0;  // 32'hfb5efeaa;
    ram_cell[      97] = 32'h0;  // 32'h6fbc9834;
    ram_cell[      98] = 32'h0;  // 32'h024ad838;
    ram_cell[      99] = 32'h0;  // 32'h14d00ce2;
    ram_cell[     100] = 32'h0;  // 32'h5cedb36e;
    ram_cell[     101] = 32'h0;  // 32'h94e17e55;
    ram_cell[     102] = 32'h0;  // 32'h9577c647;
    ram_cell[     103] = 32'h0;  // 32'h74c2a3ea;
    ram_cell[     104] = 32'h0;  // 32'h35b8a135;
    ram_cell[     105] = 32'h0;  // 32'h66cd68ec;
    ram_cell[     106] = 32'h0;  // 32'h0af87dd2;
    ram_cell[     107] = 32'h0;  // 32'hcc175b9d;
    ram_cell[     108] = 32'h0;  // 32'h5b3951c7;
    ram_cell[     109] = 32'h0;  // 32'hc3f71425;
    ram_cell[     110] = 32'h0;  // 32'h33e3a3e9;
    ram_cell[     111] = 32'h0;  // 32'h04e262c8;
    ram_cell[     112] = 32'h0;  // 32'hfd682b66;
    ram_cell[     113] = 32'h0;  // 32'h569dacde;
    ram_cell[     114] = 32'h0;  // 32'h4e59030b;
    ram_cell[     115] = 32'h0;  // 32'hae51b9b9;
    ram_cell[     116] = 32'h0;  // 32'hc9350c93;
    ram_cell[     117] = 32'h0;  // 32'h35b65ee7;
    ram_cell[     118] = 32'h0;  // 32'h289f2369;
    ram_cell[     119] = 32'h0;  // 32'h254de9d2;
    ram_cell[     120] = 32'h0;  // 32'hbc9c5bf2;
    ram_cell[     121] = 32'h0;  // 32'h61a5320c;
    ram_cell[     122] = 32'h0;  // 32'hdf1dc196;
    ram_cell[     123] = 32'h0;  // 32'h9df34314;
    ram_cell[     124] = 32'h0;  // 32'h5a4766ae;
    ram_cell[     125] = 32'h0;  // 32'h2d651b2f;
    ram_cell[     126] = 32'h0;  // 32'ha6c30774;
    ram_cell[     127] = 32'h0;  // 32'hcc3106d5;
    ram_cell[     128] = 32'h0;  // 32'h0fff554d;
    ram_cell[     129] = 32'h0;  // 32'hd2947c43;
    ram_cell[     130] = 32'h0;  // 32'hb86f2ccf;
    ram_cell[     131] = 32'h0;  // 32'h0b2c509a;
    ram_cell[     132] = 32'h0;  // 32'h64bbc77e;
    ram_cell[     133] = 32'h0;  // 32'h691ee3be;
    ram_cell[     134] = 32'h0;  // 32'h04f89291;
    ram_cell[     135] = 32'h0;  // 32'h432fc006;
    ram_cell[     136] = 32'h0;  // 32'h0fa1e4c1;
    ram_cell[     137] = 32'h0;  // 32'h462406a4;
    ram_cell[     138] = 32'h0;  // 32'hf0bf0a5c;
    ram_cell[     139] = 32'h0;  // 32'h9dbab406;
    ram_cell[     140] = 32'h0;  // 32'hd6bde9c7;
    ram_cell[     141] = 32'h0;  // 32'hae918f7a;
    ram_cell[     142] = 32'h0;  // 32'hc9603a82;
    ram_cell[     143] = 32'h0;  // 32'h9f2647e0;
    ram_cell[     144] = 32'h0;  // 32'hc4da9f4f;
    ram_cell[     145] = 32'h0;  // 32'hae306737;
    ram_cell[     146] = 32'h0;  // 32'h3bb13abb;
    ram_cell[     147] = 32'h0;  // 32'h4b976c98;
    ram_cell[     148] = 32'h0;  // 32'h7b9b05d2;
    ram_cell[     149] = 32'h0;  // 32'h75e0111d;
    ram_cell[     150] = 32'h0;  // 32'h0cfb3e43;
    ram_cell[     151] = 32'h0;  // 32'h5f120c58;
    ram_cell[     152] = 32'h0;  // 32'hf9eb64fc;
    ram_cell[     153] = 32'h0;  // 32'h084bc9f1;
    ram_cell[     154] = 32'h0;  // 32'haa7cbe6b;
    ram_cell[     155] = 32'h0;  // 32'heeb8ba14;
    ram_cell[     156] = 32'h0;  // 32'h1fad6cd0;
    ram_cell[     157] = 32'h0;  // 32'h06f1e9ae;
    ram_cell[     158] = 32'h0;  // 32'h41417ef4;
    ram_cell[     159] = 32'h0;  // 32'h75a17d27;
    ram_cell[     160] = 32'h0;  // 32'h7500e06b;
    ram_cell[     161] = 32'h0;  // 32'h127d15bd;
    ram_cell[     162] = 32'h0;  // 32'h20969d0f;
    ram_cell[     163] = 32'h0;  // 32'h21cfb3fb;
    ram_cell[     164] = 32'h0;  // 32'h067b0a89;
    ram_cell[     165] = 32'h0;  // 32'h7e5630e2;
    ram_cell[     166] = 32'h0;  // 32'h166a6fc9;
    ram_cell[     167] = 32'h0;  // 32'h0a34fcc9;
    ram_cell[     168] = 32'h0;  // 32'hd1dbbc09;
    ram_cell[     169] = 32'h0;  // 32'h160879fa;
    ram_cell[     170] = 32'h0;  // 32'h25ce825b;
    ram_cell[     171] = 32'h0;  // 32'hc234476b;
    ram_cell[     172] = 32'h0;  // 32'hc82a3b99;
    ram_cell[     173] = 32'h0;  // 32'h73b41120;
    ram_cell[     174] = 32'h0;  // 32'h4ef163de;
    ram_cell[     175] = 32'h0;  // 32'h461dee1b;
    ram_cell[     176] = 32'h0;  // 32'hcdda26bc;
    ram_cell[     177] = 32'h0;  // 32'he1c22dc9;
    ram_cell[     178] = 32'h0;  // 32'h55751381;
    ram_cell[     179] = 32'h0;  // 32'h0fcaea31;
    ram_cell[     180] = 32'h0;  // 32'h1d1bf3e0;
    ram_cell[     181] = 32'h0;  // 32'h46e5ed52;
    ram_cell[     182] = 32'h0;  // 32'hf7821a08;
    ram_cell[     183] = 32'h0;  // 32'h342927d2;
    ram_cell[     184] = 32'h0;  // 32'h34847fd8;
    ram_cell[     185] = 32'h0;  // 32'h1e31dd0e;
    ram_cell[     186] = 32'h0;  // 32'hb17e0b25;
    ram_cell[     187] = 32'h0;  // 32'h0104ea93;
    ram_cell[     188] = 32'h0;  // 32'h5e9fc4e7;
    ram_cell[     189] = 32'h0;  // 32'he0d9ee2c;
    ram_cell[     190] = 32'h0;  // 32'h81f9993b;
    ram_cell[     191] = 32'h0;  // 32'h7d127ed6;
    ram_cell[     192] = 32'h0;  // 32'ha700f86f;
    ram_cell[     193] = 32'h0;  // 32'h77b8bc82;
    ram_cell[     194] = 32'h0;  // 32'h33c67dd7;
    ram_cell[     195] = 32'h0;  // 32'h7eda8561;
    ram_cell[     196] = 32'h0;  // 32'h12f43ff1;
    ram_cell[     197] = 32'h0;  // 32'hacf9081a;
    ram_cell[     198] = 32'h0;  // 32'h6affa00e;
    ram_cell[     199] = 32'h0;  // 32'h51a1a2c9;
    ram_cell[     200] = 32'h0;  // 32'h046c3f06;
    ram_cell[     201] = 32'h0;  // 32'hbfc0bddc;
    ram_cell[     202] = 32'h0;  // 32'hb6e26f7c;
    ram_cell[     203] = 32'h0;  // 32'h56cd1fa8;
    ram_cell[     204] = 32'h0;  // 32'heed73470;
    ram_cell[     205] = 32'h0;  // 32'h56e8d9cd;
    ram_cell[     206] = 32'h0;  // 32'h089f5f97;
    ram_cell[     207] = 32'h0;  // 32'h778bcef2;
    ram_cell[     208] = 32'h0;  // 32'h70d1d450;
    ram_cell[     209] = 32'h0;  // 32'h549be943;
    ram_cell[     210] = 32'h0;  // 32'h2c75907f;
    ram_cell[     211] = 32'h0;  // 32'hdfc4b897;
    ram_cell[     212] = 32'h0;  // 32'h574cb3b5;
    ram_cell[     213] = 32'h0;  // 32'h8635014f;
    ram_cell[     214] = 32'h0;  // 32'h953d587f;
    ram_cell[     215] = 32'h0;  // 32'ha7ccc9b1;
    ram_cell[     216] = 32'h0;  // 32'h59dfd13d;
    ram_cell[     217] = 32'h0;  // 32'hac4657b8;
    ram_cell[     218] = 32'h0;  // 32'hd48fdc41;
    ram_cell[     219] = 32'h0;  // 32'h4169db8d;
    ram_cell[     220] = 32'h0;  // 32'h64e35a90;
    ram_cell[     221] = 32'h0;  // 32'hfb9343ff;
    ram_cell[     222] = 32'h0;  // 32'hc3d49358;
    ram_cell[     223] = 32'h0;  // 32'h5c4c00c2;
    ram_cell[     224] = 32'h0;  // 32'h77b17be0;
    ram_cell[     225] = 32'h0;  // 32'h80624802;
    ram_cell[     226] = 32'h0;  // 32'hfc1c6c6b;
    ram_cell[     227] = 32'h0;  // 32'h202e9bd7;
    ram_cell[     228] = 32'h0;  // 32'ha68ee21c;
    ram_cell[     229] = 32'h0;  // 32'h57d7635c;
    ram_cell[     230] = 32'h0;  // 32'h2a3e2ceb;
    ram_cell[     231] = 32'h0;  // 32'h18861fba;
    ram_cell[     232] = 32'h0;  // 32'he9f88b6e;
    ram_cell[     233] = 32'h0;  // 32'h55275388;
    ram_cell[     234] = 32'h0;  // 32'h473e48bb;
    ram_cell[     235] = 32'h0;  // 32'h8df53027;
    ram_cell[     236] = 32'h0;  // 32'h255b682b;
    ram_cell[     237] = 32'h0;  // 32'h8cfc85a8;
    ram_cell[     238] = 32'h0;  // 32'hf829d29d;
    ram_cell[     239] = 32'h0;  // 32'heaa8cd68;
    ram_cell[     240] = 32'h0;  // 32'he958232e;
    ram_cell[     241] = 32'h0;  // 32'hadc314ab;
    ram_cell[     242] = 32'h0;  // 32'h397f4267;
    ram_cell[     243] = 32'h0;  // 32'hdf071b26;
    ram_cell[     244] = 32'h0;  // 32'hd6ef1f79;
    ram_cell[     245] = 32'h0;  // 32'h4c3fc4e7;
    ram_cell[     246] = 32'h0;  // 32'hba630722;
    ram_cell[     247] = 32'h0;  // 32'h61af984c;
    ram_cell[     248] = 32'h0;  // 32'h25605b70;
    ram_cell[     249] = 32'h0;  // 32'h76a81db4;
    ram_cell[     250] = 32'h0;  // 32'hee65af5b;
    ram_cell[     251] = 32'h0;  // 32'h8c4f7a5c;
    ram_cell[     252] = 32'h0;  // 32'hc21c1ccb;
    ram_cell[     253] = 32'h0;  // 32'h2a775452;
    ram_cell[     254] = 32'h0;  // 32'hc50e7d6a;
    ram_cell[     255] = 32'h0;  // 32'h8ad7b207;
    // src matrix A
    ram_cell[     256] = 32'h25289341;
    ram_cell[     257] = 32'h32c12c25;
    ram_cell[     258] = 32'hae76943a;
    ram_cell[     259] = 32'h859bf6aa;
    ram_cell[     260] = 32'h63392035;
    ram_cell[     261] = 32'he3e9dc8c;
    ram_cell[     262] = 32'hb63561f7;
    ram_cell[     263] = 32'hde7a161e;
    ram_cell[     264] = 32'h8c9087f2;
    ram_cell[     265] = 32'hb8dcf9ff;
    ram_cell[     266] = 32'h5c1e5eac;
    ram_cell[     267] = 32'h7d5370a4;
    ram_cell[     268] = 32'hb0fb013a;
    ram_cell[     269] = 32'h083af099;
    ram_cell[     270] = 32'h109b7a10;
    ram_cell[     271] = 32'h8bbaa745;
    ram_cell[     272] = 32'he9c3230f;
    ram_cell[     273] = 32'h94de907b;
    ram_cell[     274] = 32'heae2135f;
    ram_cell[     275] = 32'hec58777d;
    ram_cell[     276] = 32'h5a09062d;
    ram_cell[     277] = 32'hf92bbdfa;
    ram_cell[     278] = 32'hd1646776;
    ram_cell[     279] = 32'he59a460a;
    ram_cell[     280] = 32'h3ba4f9e3;
    ram_cell[     281] = 32'h99d230f1;
    ram_cell[     282] = 32'h612e4fd0;
    ram_cell[     283] = 32'h7c84ba07;
    ram_cell[     284] = 32'h52ef1181;
    ram_cell[     285] = 32'h23ca8918;
    ram_cell[     286] = 32'h0deeaf4c;
    ram_cell[     287] = 32'hd57a5b2d;
    ram_cell[     288] = 32'hc4415cb0;
    ram_cell[     289] = 32'h3212cb35;
    ram_cell[     290] = 32'hd730d0f6;
    ram_cell[     291] = 32'h5fc9682b;
    ram_cell[     292] = 32'hbc7366e9;
    ram_cell[     293] = 32'hf08acf73;
    ram_cell[     294] = 32'h8f670f69;
    ram_cell[     295] = 32'h46615b1b;
    ram_cell[     296] = 32'h264c5781;
    ram_cell[     297] = 32'h4ef7c098;
    ram_cell[     298] = 32'h32b75be6;
    ram_cell[     299] = 32'he72ddb0a;
    ram_cell[     300] = 32'h16e6ab93;
    ram_cell[     301] = 32'h8c4a9ab4;
    ram_cell[     302] = 32'h8743753d;
    ram_cell[     303] = 32'h4183b328;
    ram_cell[     304] = 32'h28931412;
    ram_cell[     305] = 32'h15fc4f55;
    ram_cell[     306] = 32'h7e96f388;
    ram_cell[     307] = 32'ha310503b;
    ram_cell[     308] = 32'h10a4dbf3;
    ram_cell[     309] = 32'hfa310fe0;
    ram_cell[     310] = 32'h0b87d783;
    ram_cell[     311] = 32'hecd44232;
    ram_cell[     312] = 32'h6003d3cc;
    ram_cell[     313] = 32'h0775e722;
    ram_cell[     314] = 32'hf4ec95ad;
    ram_cell[     315] = 32'h3f3e3c25;
    ram_cell[     316] = 32'hbdd8bafc;
    ram_cell[     317] = 32'hab153f0e;
    ram_cell[     318] = 32'h2acd302d;
    ram_cell[     319] = 32'hb74c6af4;
    ram_cell[     320] = 32'h043fac99;
    ram_cell[     321] = 32'hbb89d84b;
    ram_cell[     322] = 32'h756079af;
    ram_cell[     323] = 32'hf6d1a16d;
    ram_cell[     324] = 32'hff64ee5c;
    ram_cell[     325] = 32'hd743248e;
    ram_cell[     326] = 32'h6eeb2129;
    ram_cell[     327] = 32'h7546c44e;
    ram_cell[     328] = 32'h40b02ada;
    ram_cell[     329] = 32'h533babc9;
    ram_cell[     330] = 32'h515ec375;
    ram_cell[     331] = 32'h5e83f209;
    ram_cell[     332] = 32'h4edcde89;
    ram_cell[     333] = 32'hb251dbe7;
    ram_cell[     334] = 32'h48285901;
    ram_cell[     335] = 32'h8d254b60;
    ram_cell[     336] = 32'hf53de831;
    ram_cell[     337] = 32'h7640a146;
    ram_cell[     338] = 32'h959ac476;
    ram_cell[     339] = 32'hac86ef8f;
    ram_cell[     340] = 32'hb1c49845;
    ram_cell[     341] = 32'h8de581c0;
    ram_cell[     342] = 32'h95d3811a;
    ram_cell[     343] = 32'h4ef11efb;
    ram_cell[     344] = 32'h174f2154;
    ram_cell[     345] = 32'hca1c1ed5;
    ram_cell[     346] = 32'h6f286681;
    ram_cell[     347] = 32'h954229a7;
    ram_cell[     348] = 32'h541a37dd;
    ram_cell[     349] = 32'h27e0d9ad;
    ram_cell[     350] = 32'hacfe525b;
    ram_cell[     351] = 32'h59f52778;
    ram_cell[     352] = 32'ha7f1caf9;
    ram_cell[     353] = 32'h367b3cff;
    ram_cell[     354] = 32'h3c02efaf;
    ram_cell[     355] = 32'ha9b8b1b8;
    ram_cell[     356] = 32'hb9961074;
    ram_cell[     357] = 32'h2b966ba0;
    ram_cell[     358] = 32'h0a85acae;
    ram_cell[     359] = 32'h704c246e;
    ram_cell[     360] = 32'h3fe7bd01;
    ram_cell[     361] = 32'h22ce038e;
    ram_cell[     362] = 32'h4c6a633c;
    ram_cell[     363] = 32'h7fd6e189;
    ram_cell[     364] = 32'hc4ba97d4;
    ram_cell[     365] = 32'ha3a31902;
    ram_cell[     366] = 32'h390aa76b;
    ram_cell[     367] = 32'h827b9c9b;
    ram_cell[     368] = 32'h0d9bc239;
    ram_cell[     369] = 32'ha196f237;
    ram_cell[     370] = 32'h83d5ca6b;
    ram_cell[     371] = 32'h04a93ef1;
    ram_cell[     372] = 32'h080a6f5c;
    ram_cell[     373] = 32'hb6e9d6ad;
    ram_cell[     374] = 32'h10ef4fc1;
    ram_cell[     375] = 32'h8b1ca76e;
    ram_cell[     376] = 32'h1b04ac55;
    ram_cell[     377] = 32'h14108d83;
    ram_cell[     378] = 32'hdbb20ac2;
    ram_cell[     379] = 32'h739e416d;
    ram_cell[     380] = 32'haf3dad6a;
    ram_cell[     381] = 32'he713ee91;
    ram_cell[     382] = 32'h92e489f1;
    ram_cell[     383] = 32'h2c639bf0;
    ram_cell[     384] = 32'hd6887ce1;
    ram_cell[     385] = 32'h6e068ef7;
    ram_cell[     386] = 32'hd8f43de6;
    ram_cell[     387] = 32'hc11618aa;
    ram_cell[     388] = 32'h1864bbf3;
    ram_cell[     389] = 32'hdbea319f;
    ram_cell[     390] = 32'hefdf381e;
    ram_cell[     391] = 32'hf7b89f74;
    ram_cell[     392] = 32'h1801ebf4;
    ram_cell[     393] = 32'hc0edb8bc;
    ram_cell[     394] = 32'hd0852008;
    ram_cell[     395] = 32'h88cf804d;
    ram_cell[     396] = 32'hd8a65f8f;
    ram_cell[     397] = 32'h30975244;
    ram_cell[     398] = 32'hc265d023;
    ram_cell[     399] = 32'h1142ee11;
    ram_cell[     400] = 32'h58210f0f;
    ram_cell[     401] = 32'h6a811188;
    ram_cell[     402] = 32'h80cc92f3;
    ram_cell[     403] = 32'hcbbdeeb4;
    ram_cell[     404] = 32'h641de3f2;
    ram_cell[     405] = 32'h1933679a;
    ram_cell[     406] = 32'h40372d1a;
    ram_cell[     407] = 32'h967c076e;
    ram_cell[     408] = 32'hcf4bcc53;
    ram_cell[     409] = 32'h208fd044;
    ram_cell[     410] = 32'h4241c40d;
    ram_cell[     411] = 32'h0cbccc70;
    ram_cell[     412] = 32'h69e70591;
    ram_cell[     413] = 32'h606a1e57;
    ram_cell[     414] = 32'h5ba1c8f2;
    ram_cell[     415] = 32'ha5314bfc;
    ram_cell[     416] = 32'h14d4480c;
    ram_cell[     417] = 32'h16236ca2;
    ram_cell[     418] = 32'hb523bd8d;
    ram_cell[     419] = 32'h80e53b81;
    ram_cell[     420] = 32'h432a11f3;
    ram_cell[     421] = 32'h94c463be;
    ram_cell[     422] = 32'h0ff2e896;
    ram_cell[     423] = 32'h81a14337;
    ram_cell[     424] = 32'hfa559b84;
    ram_cell[     425] = 32'hec616a1b;
    ram_cell[     426] = 32'h8815af4c;
    ram_cell[     427] = 32'h6b581d7c;
    ram_cell[     428] = 32'h2520a197;
    ram_cell[     429] = 32'h7b080933;
    ram_cell[     430] = 32'hefb69d40;
    ram_cell[     431] = 32'hba245638;
    ram_cell[     432] = 32'h3ada7d63;
    ram_cell[     433] = 32'h11486d79;
    ram_cell[     434] = 32'hb9a0344f;
    ram_cell[     435] = 32'h417b2d8e;
    ram_cell[     436] = 32'h4482599d;
    ram_cell[     437] = 32'hff39fec3;
    ram_cell[     438] = 32'hbae76faa;
    ram_cell[     439] = 32'h719c1cab;
    ram_cell[     440] = 32'he3f50ef5;
    ram_cell[     441] = 32'hee9cd63f;
    ram_cell[     442] = 32'h51c99d1a;
    ram_cell[     443] = 32'h1bfaeb14;
    ram_cell[     444] = 32'h32f0d686;
    ram_cell[     445] = 32'h2d796d2c;
    ram_cell[     446] = 32'h8dd101fc;
    ram_cell[     447] = 32'h02b234dc;
    ram_cell[     448] = 32'hd0980803;
    ram_cell[     449] = 32'h420e782c;
    ram_cell[     450] = 32'hbd40e729;
    ram_cell[     451] = 32'h45a04012;
    ram_cell[     452] = 32'h24602fcf;
    ram_cell[     453] = 32'h546f9d0c;
    ram_cell[     454] = 32'hb033dd8a;
    ram_cell[     455] = 32'h5cdf363d;
    ram_cell[     456] = 32'h1e82a544;
    ram_cell[     457] = 32'h76060cc5;
    ram_cell[     458] = 32'hab259bbf;
    ram_cell[     459] = 32'h8cbedeab;
    ram_cell[     460] = 32'ha3e1885e;
    ram_cell[     461] = 32'h12030133;
    ram_cell[     462] = 32'h956c43aa;
    ram_cell[     463] = 32'hdb391c2d;
    ram_cell[     464] = 32'h0e1592c5;
    ram_cell[     465] = 32'h40fbe7af;
    ram_cell[     466] = 32'h4c53df06;
    ram_cell[     467] = 32'h4f4932c0;
    ram_cell[     468] = 32'h8c1ef358;
    ram_cell[     469] = 32'hc85119e5;
    ram_cell[     470] = 32'h7bcbb734;
    ram_cell[     471] = 32'h750dd86e;
    ram_cell[     472] = 32'hff83cd9b;
    ram_cell[     473] = 32'h98f7e026;
    ram_cell[     474] = 32'h9d8b325b;
    ram_cell[     475] = 32'haa422ba6;
    ram_cell[     476] = 32'h9b0f2809;
    ram_cell[     477] = 32'h31ca07ad;
    ram_cell[     478] = 32'hfae384ee;
    ram_cell[     479] = 32'hfdbbca24;
    ram_cell[     480] = 32'h3e86abc3;
    ram_cell[     481] = 32'hadbfbc84;
    ram_cell[     482] = 32'h2c2d7d35;
    ram_cell[     483] = 32'h8738abc3;
    ram_cell[     484] = 32'h4649d741;
    ram_cell[     485] = 32'hb8cafc8c;
    ram_cell[     486] = 32'h68f4bf82;
    ram_cell[     487] = 32'hc54835c7;
    ram_cell[     488] = 32'heb1c39b2;
    ram_cell[     489] = 32'hf99b2085;
    ram_cell[     490] = 32'hc7d57995;
    ram_cell[     491] = 32'h0a9ada27;
    ram_cell[     492] = 32'h502c5567;
    ram_cell[     493] = 32'h1b250238;
    ram_cell[     494] = 32'hd506f19d;
    ram_cell[     495] = 32'h211921f0;
    ram_cell[     496] = 32'h5c426f95;
    ram_cell[     497] = 32'hbb8ca265;
    ram_cell[     498] = 32'hdd0e4ed7;
    ram_cell[     499] = 32'hebb1f60c;
    ram_cell[     500] = 32'ha52a6b00;
    ram_cell[     501] = 32'hfc8ce4dd;
    ram_cell[     502] = 32'hdaf16dc1;
    ram_cell[     503] = 32'hc597e354;
    ram_cell[     504] = 32'hbe03c055;
    ram_cell[     505] = 32'hff654212;
    ram_cell[     506] = 32'h35d3fc33;
    ram_cell[     507] = 32'h3f8c4369;
    ram_cell[     508] = 32'hf0a1a1be;
    ram_cell[     509] = 32'h836dd8e9;
    ram_cell[     510] = 32'he9f00ebf;
    ram_cell[     511] = 32'h7ca266b9;
    // src matrix B
    ram_cell[     512] = 32'he8935bdb;
    ram_cell[     513] = 32'h48a06609;
    ram_cell[     514] = 32'hbfde9bec;
    ram_cell[     515] = 32'h54e150c6;
    ram_cell[     516] = 32'hae5834a8;
    ram_cell[     517] = 32'hb4f429eb;
    ram_cell[     518] = 32'hb009d94e;
    ram_cell[     519] = 32'h4ad6c232;
    ram_cell[     520] = 32'h1a26ae83;
    ram_cell[     521] = 32'hbf422f50;
    ram_cell[     522] = 32'h2fc041aa;
    ram_cell[     523] = 32'hb2b1f639;
    ram_cell[     524] = 32'h0c170d30;
    ram_cell[     525] = 32'h59988cd7;
    ram_cell[     526] = 32'h2310df45;
    ram_cell[     527] = 32'h7fd475ae;
    ram_cell[     528] = 32'h27ad17b8;
    ram_cell[     529] = 32'hc68e99e9;
    ram_cell[     530] = 32'hc34876fb;
    ram_cell[     531] = 32'hbcf6c020;
    ram_cell[     532] = 32'hd1a2d744;
    ram_cell[     533] = 32'he8d4235a;
    ram_cell[     534] = 32'h4aef1e59;
    ram_cell[     535] = 32'h1c650e69;
    ram_cell[     536] = 32'h8bdab9c8;
    ram_cell[     537] = 32'hb8557e5a;
    ram_cell[     538] = 32'h06455739;
    ram_cell[     539] = 32'h04d8fe98;
    ram_cell[     540] = 32'h28d83d66;
    ram_cell[     541] = 32'h2cbefa03;
    ram_cell[     542] = 32'h7ce50418;
    ram_cell[     543] = 32'ha2a18b24;
    ram_cell[     544] = 32'h5e1fc5c9;
    ram_cell[     545] = 32'h26469762;
    ram_cell[     546] = 32'h28a0bc35;
    ram_cell[     547] = 32'h050db0e3;
    ram_cell[     548] = 32'h02769a00;
    ram_cell[     549] = 32'hba03d374;
    ram_cell[     550] = 32'h552c7c59;
    ram_cell[     551] = 32'h71b21624;
    ram_cell[     552] = 32'hf55282a4;
    ram_cell[     553] = 32'heb592586;
    ram_cell[     554] = 32'h8dc0b8ad;
    ram_cell[     555] = 32'ha72b567d;
    ram_cell[     556] = 32'hb584e020;
    ram_cell[     557] = 32'he7fa5c9b;
    ram_cell[     558] = 32'h4d05932e;
    ram_cell[     559] = 32'h7969e9ee;
    ram_cell[     560] = 32'he8ab22c0;
    ram_cell[     561] = 32'ha66d7ca3;
    ram_cell[     562] = 32'hdfbc276b;
    ram_cell[     563] = 32'h05f111d5;
    ram_cell[     564] = 32'h15364e19;
    ram_cell[     565] = 32'hf3c2f94f;
    ram_cell[     566] = 32'h5a8f5cb8;
    ram_cell[     567] = 32'h39b811ef;
    ram_cell[     568] = 32'hb3cb6b09;
    ram_cell[     569] = 32'h77e84be9;
    ram_cell[     570] = 32'hb0ed77c8;
    ram_cell[     571] = 32'h190cd121;
    ram_cell[     572] = 32'h5bece9c4;
    ram_cell[     573] = 32'h2ee4767e;
    ram_cell[     574] = 32'h632a41f4;
    ram_cell[     575] = 32'h3c79a36c;
    ram_cell[     576] = 32'hd045fe18;
    ram_cell[     577] = 32'h51bcab6d;
    ram_cell[     578] = 32'hb24126f0;
    ram_cell[     579] = 32'h8cc3a499;
    ram_cell[     580] = 32'h4b1f2990;
    ram_cell[     581] = 32'h61eeac27;
    ram_cell[     582] = 32'h2392ff3d;
    ram_cell[     583] = 32'h5f437508;
    ram_cell[     584] = 32'hb8cd0bca;
    ram_cell[     585] = 32'h9eb30f5f;
    ram_cell[     586] = 32'hef5ac318;
    ram_cell[     587] = 32'hc7e5c7a1;
    ram_cell[     588] = 32'h2fd640c5;
    ram_cell[     589] = 32'h73a282a8;
    ram_cell[     590] = 32'h002ace75;
    ram_cell[     591] = 32'h8a6399a9;
    ram_cell[     592] = 32'h5d27d92a;
    ram_cell[     593] = 32'h6139f967;
    ram_cell[     594] = 32'h8fd65078;
    ram_cell[     595] = 32'h446fc7a2;
    ram_cell[     596] = 32'h2d486e49;
    ram_cell[     597] = 32'h0bdca56e;
    ram_cell[     598] = 32'hd030f856;
    ram_cell[     599] = 32'h0ddb04f6;
    ram_cell[     600] = 32'h76237c77;
    ram_cell[     601] = 32'h8213c573;
    ram_cell[     602] = 32'h30eb9640;
    ram_cell[     603] = 32'hb229bb4a;
    ram_cell[     604] = 32'h6972bb36;
    ram_cell[     605] = 32'h63ba9e9b;
    ram_cell[     606] = 32'h0e593186;
    ram_cell[     607] = 32'hc5b68299;
    ram_cell[     608] = 32'h34ed39cd;
    ram_cell[     609] = 32'h40a74f63;
    ram_cell[     610] = 32'hd2a4724b;
    ram_cell[     611] = 32'h06cbe6b3;
    ram_cell[     612] = 32'h3621355d;
    ram_cell[     613] = 32'h416e6248;
    ram_cell[     614] = 32'h6f824e2f;
    ram_cell[     615] = 32'ha2fa0e94;
    ram_cell[     616] = 32'h5ab44092;
    ram_cell[     617] = 32'h32dbeb82;
    ram_cell[     618] = 32'hd85b13c6;
    ram_cell[     619] = 32'h1c887728;
    ram_cell[     620] = 32'hdd295d8b;
    ram_cell[     621] = 32'h4feb891b;
    ram_cell[     622] = 32'h574011d8;
    ram_cell[     623] = 32'hc85782c3;
    ram_cell[     624] = 32'hb93526d8;
    ram_cell[     625] = 32'h7fe19bb6;
    ram_cell[     626] = 32'h63b8ca74;
    ram_cell[     627] = 32'h7c02faf5;
    ram_cell[     628] = 32'h7aeba68b;
    ram_cell[     629] = 32'h42029ece;
    ram_cell[     630] = 32'hfe8955f5;
    ram_cell[     631] = 32'h310e3189;
    ram_cell[     632] = 32'h689f2de4;
    ram_cell[     633] = 32'h056ecc8b;
    ram_cell[     634] = 32'h9bf592e2;
    ram_cell[     635] = 32'h76cfc9d6;
    ram_cell[     636] = 32'h96cb3b77;
    ram_cell[     637] = 32'hb0281b58;
    ram_cell[     638] = 32'h462ba449;
    ram_cell[     639] = 32'hf90c1d4b;
    ram_cell[     640] = 32'h5b305ff7;
    ram_cell[     641] = 32'h98cb8bc5;
    ram_cell[     642] = 32'h3c0816f7;
    ram_cell[     643] = 32'h27aefeb9;
    ram_cell[     644] = 32'h0c5dc1fa;
    ram_cell[     645] = 32'h4fd4cdf3;
    ram_cell[     646] = 32'h32f6e21e;
    ram_cell[     647] = 32'h8c3ec2d4;
    ram_cell[     648] = 32'h442d495f;
    ram_cell[     649] = 32'h1c2f54d2;
    ram_cell[     650] = 32'h51da4f19;
    ram_cell[     651] = 32'h77d81d91;
    ram_cell[     652] = 32'h43b78924;
    ram_cell[     653] = 32'hc8502a8d;
    ram_cell[     654] = 32'hd8e3dca9;
    ram_cell[     655] = 32'hb0aadf26;
    ram_cell[     656] = 32'ha7243b77;
    ram_cell[     657] = 32'hc8294e0a;
    ram_cell[     658] = 32'h9eb2ca14;
    ram_cell[     659] = 32'h9adb7d65;
    ram_cell[     660] = 32'h0a6241aa;
    ram_cell[     661] = 32'hea9fa865;
    ram_cell[     662] = 32'hdd47556a;
    ram_cell[     663] = 32'h403e74c6;
    ram_cell[     664] = 32'h9ccd48a1;
    ram_cell[     665] = 32'hc156094f;
    ram_cell[     666] = 32'h6be16890;
    ram_cell[     667] = 32'hf35dea93;
    ram_cell[     668] = 32'h3b8c876b;
    ram_cell[     669] = 32'h77d178b7;
    ram_cell[     670] = 32'hc99d4a33;
    ram_cell[     671] = 32'hd2cfe827;
    ram_cell[     672] = 32'hb6d093db;
    ram_cell[     673] = 32'hef5f0dc2;
    ram_cell[     674] = 32'h67aba764;
    ram_cell[     675] = 32'hdd1da2d6;
    ram_cell[     676] = 32'h1ba7fc35;
    ram_cell[     677] = 32'h173767be;
    ram_cell[     678] = 32'h8f2ed04a;
    ram_cell[     679] = 32'h46bf8daf;
    ram_cell[     680] = 32'hde05059f;
    ram_cell[     681] = 32'h33796857;
    ram_cell[     682] = 32'h4aa5d7bf;
    ram_cell[     683] = 32'h16642b7c;
    ram_cell[     684] = 32'h5fcd5a7c;
    ram_cell[     685] = 32'hddb063df;
    ram_cell[     686] = 32'hc9c23c51;
    ram_cell[     687] = 32'h3ac46ea7;
    ram_cell[     688] = 32'hb00f37bb;
    ram_cell[     689] = 32'h09b6abd7;
    ram_cell[     690] = 32'h931404d3;
    ram_cell[     691] = 32'he8dd0833;
    ram_cell[     692] = 32'hcb67edf5;
    ram_cell[     693] = 32'h5aa42353;
    ram_cell[     694] = 32'h01dbd818;
    ram_cell[     695] = 32'he4884638;
    ram_cell[     696] = 32'h17f10ab7;
    ram_cell[     697] = 32'h801855a3;
    ram_cell[     698] = 32'h6bfb790c;
    ram_cell[     699] = 32'h6b092e1f;
    ram_cell[     700] = 32'hc54f4b4a;
    ram_cell[     701] = 32'h1df9f146;
    ram_cell[     702] = 32'hc077a576;
    ram_cell[     703] = 32'he5975fda;
    ram_cell[     704] = 32'h39ac358d;
    ram_cell[     705] = 32'h1053dd8a;
    ram_cell[     706] = 32'hcba903cb;
    ram_cell[     707] = 32'he981d4b3;
    ram_cell[     708] = 32'h97c6c3cf;
    ram_cell[     709] = 32'h76c3432d;
    ram_cell[     710] = 32'hc21d9e62;
    ram_cell[     711] = 32'hf4a8b4ce;
    ram_cell[     712] = 32'h3e48c3b0;
    ram_cell[     713] = 32'hf1eb5cda;
    ram_cell[     714] = 32'hfa7bff7e;
    ram_cell[     715] = 32'h6a1e36f0;
    ram_cell[     716] = 32'hc57ae7c9;
    ram_cell[     717] = 32'h0bacebbc;
    ram_cell[     718] = 32'ha7f12305;
    ram_cell[     719] = 32'h2f57ba22;
    ram_cell[     720] = 32'h0f0fbb50;
    ram_cell[     721] = 32'h82bf18b5;
    ram_cell[     722] = 32'he1a60c6a;
    ram_cell[     723] = 32'hd29e92d7;
    ram_cell[     724] = 32'h4c342050;
    ram_cell[     725] = 32'h40c22526;
    ram_cell[     726] = 32'hdc1f470a;
    ram_cell[     727] = 32'h1a02f51d;
    ram_cell[     728] = 32'h14c804a1;
    ram_cell[     729] = 32'hb2dcbb34;
    ram_cell[     730] = 32'h7fc5021c;
    ram_cell[     731] = 32'h7a5e5eb5;
    ram_cell[     732] = 32'h195f988f;
    ram_cell[     733] = 32'h2a495c6e;
    ram_cell[     734] = 32'hee2f759a;
    ram_cell[     735] = 32'hafd0bf28;
    ram_cell[     736] = 32'h357957f4;
    ram_cell[     737] = 32'h109aac38;
    ram_cell[     738] = 32'h14e7780f;
    ram_cell[     739] = 32'h3a25ddee;
    ram_cell[     740] = 32'hd8bfce39;
    ram_cell[     741] = 32'h7302dd6e;
    ram_cell[     742] = 32'h7be99f50;
    ram_cell[     743] = 32'hf73a48c7;
    ram_cell[     744] = 32'h2f740e4f;
    ram_cell[     745] = 32'h6e3f240c;
    ram_cell[     746] = 32'hc6371aab;
    ram_cell[     747] = 32'h3090a8d5;
    ram_cell[     748] = 32'h93eac4bb;
    ram_cell[     749] = 32'hca783fcc;
    ram_cell[     750] = 32'h985c1a5f;
    ram_cell[     751] = 32'hd4734c18;
    ram_cell[     752] = 32'h504cfb80;
    ram_cell[     753] = 32'h3515f1c4;
    ram_cell[     754] = 32'hb1cae4f3;
    ram_cell[     755] = 32'hb5726843;
    ram_cell[     756] = 32'h2f4f9738;
    ram_cell[     757] = 32'hf28062ba;
    ram_cell[     758] = 32'hc18a7cc3;
    ram_cell[     759] = 32'h2b277ab8;
    ram_cell[     760] = 32'hb4d35925;
    ram_cell[     761] = 32'h710c06f9;
    ram_cell[     762] = 32'hab4760e0;
    ram_cell[     763] = 32'hf02d6458;
    ram_cell[     764] = 32'h282b2326;
    ram_cell[     765] = 32'h724d765f;
    ram_cell[     766] = 32'hae4fb5ea;
    ram_cell[     767] = 32'h00b66824;
end

endmodule

